module state_transitions(
	input logic [1:0] coins,
	input logic [3:0] currentState,
	output logic [3:0] newState
);



endmodule
module main(input logic switch[2:0], buttons[1:0], realClk);

and();
endmodule
module main(
	input logic [2:0] switches, 
	input logic [1:0] buttons, 
	input logic realClk, 
	output logic [4:0] outputLED, 
	output logic [3:0] stateLED, 
	output logic [6:0] stateDisplay, changeDisplay
);


endmodule
module state3PlusTo0 (
	input logic [3:0] state,
	output lgoic [1:0] tinyState
);



endmodule